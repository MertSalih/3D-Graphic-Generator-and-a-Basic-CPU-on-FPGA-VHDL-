library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
 
entity InstReg is
    Port (order: in std_logic_vector(7 downto 0);
		  inst: out std_logic_vector(31 downto 0));
end InstReg;

architecture Behavioral of InstReg is

type reg256_32 is array  (0 to 255) of std_logic_vector(31 downto 0);
signal reg: reg256_32:=(
"11000000000000000000000000000000",
"11000000000000001000000000000001",
"11010111110000000000000010000000",
"11001000000000000000000000001001",
"10101000000100100000000000000001",
"10101000000100000000000000000000",
"11111000000000000000000000000000",
"11111000000000000000000000000000",
"11000000000000110000000000000001",
"10101000000001000000000000000000",
"10101000000001001000000000101010",
"10101000000001100000000000000001",
"10101000000001101000000000101011",
"11010111110000000000000000001000",
"11001000000000000000000000010010",
"01011001000001010000000000000001",
"01011001001001011000000000000001",
"11001000000000000000000000010110",
"11010111110000000000000000000100",
"11001000000000000000000000101111",
"01010001000001010000000000000001",
"01010001001001011000000000000001",
"10110001010000000000000000000000",
"10110001010000000000000000000110",
"10110001010000000000000000011000",
"10110001010000000000000000011110",
"10110001010000000000000000110000",
"10110001010000000000000000110110",
"10110001010000000000000000000011",
"10110001010000000000000000010101",
"10110001010000000000000000011011",
"10110001010000000000000000101101",
"10110001010000000000000000110011",
"10110001010000000000000000111001",
"10110001011000000000000000001100",
"10110001011000000000000000010010",
"10110001011000000000000000100100",
"10110001011000000000000000101010",
"10110001011000000000000000111100",
"10110001011000000000000001000010",
"10110001011000000000000000001001",
"10110001011000000000000000001111",
"10110001011000000000000000100001",
"10110001011000000000000000100111",
"10110001011000000000000000111111",
"10110001011000000000000001000101",
"11001000000000000000000001010000",
"11010111110000000000000000000010",
"11001000000000000000000000110100",
"01011001100001110000000000000001",
"01011001101001111000000000000001",
"11001000000000000000000000111000",
"11010111110000000000000000000001",
"11001000000000000000000001010000",
"01010001100001110000000000000001",
"01010001101001111000000000000001",
"10110001110000000000000000000001",
"10110001110000000000000000000111",
"10110001110000000000000000001101",
"10110001110000000000000000010011",
"10110001110000000000000000110001",
"10110001110000000000000000110111",
"10110001110000000000000000111101",
"10110001110000000000000001000011",
"10110001110000000000000000000100",
"10110001110000000000000000001010",
"10110001110000000000000000010000",
"10110001110000000000000000010110",
"10110001111000000000000000011001",
"10110001111000000000000000011111",
"10110001111000000000000000100101",
"10110001111000000000000000101011",
"10110001111000000000000000011100",
"10110001111000000000000000100010",
"10110001111000000000000000101000",
"10110001111000000000000000101110",
"10110001111000000000000000110100",
"10110001111000000000000000111010",
"10110001111000000000000001000000",
"10110001111000000000000001000110",
"10110111111000000000000010000000",
"11001000000000000000000001010111",
"10101000000100010000000001001000",
"10101000000100101000000001001001",
"11111000000000000000000000000000",
"11111000000000000000000000000000",
"11000000000000111000000000000001",
"10101000000010000000000001001000",
"10101000000010001000000001110010",
"10101000000010100000000001001001",
"10101000000010101000000001110011",
"11010111111000000000000000001000",
"11001000000000000000000001100000",
"01011010000010010000000000000001",
"01011010001010011000000000000001",
"11001000000000000000000001100100",
"11010111111000000000000000000100",
"11001000000000000000000001111101",
"01010010000010010000000000000001",
"01010010001010011000000000000001",
"10110010010000000000000001001000",
"10110010010000000000000001001110",
"10110010010000000000000001100000",
"10110010010000000000000001100110",
"10110010010000000000000001111000",
"10110010010000000000000001111110",
"10110010010000000000000001001011",
"10110010010000000000000001011101",
"10110010010000000000000001100011",
"10110010010000000000000001110101",
"10110010010000000000000001111011",
"10110010010000000000000010000001",
"10110010011000000000000001010100",
"10110010011000000000000001011010",
"10110010011000000000000001101100",
"10110010011000000000000001110010",
"10110010011000000000000010000100",
"10110010011000000000000010001010",
"10110010011000000000000001010001",
"10110010011000000000000001010111",
"10110010011000000000000001101001",
"10110010011000000000000001101111",
"10110010011000000000000010000111",
"10110010011000000000000010001101",
"11001000000000000000000010011110",
"11010111111000000000000000000010",
"11001000000000000000000010000010",
"01011010100010110000000000000001",
"01011010101010111000000000000001",
"11001000000000000000000010000110",
"11010111111000000000000000000001",
"11001000000000000000000010011110",
"01010010100010110000000000000001",
"01010010101010111000000000000001",
"10110010110000000000000001001001",
"10110010110000000000000001001111",
"10110010110000000000000001010101",
"10110010110000000000000001011011",
"10110010110000000000000001111001",
"10110010110000000000000001111111",
"10110010110000000000000010000101",
"10110010110000000000000010001011",
"10110010110000000000000001001100",
"10110010110000000000000001010010",
"10110010110000000000000001011000",
"10110010110000000000000001011110",
"10110010111000000000000001100001",
"10110010111000000000000001100111",
"10110010111000000000000001101101",
"10110010111000000000000001110011",
"10110010111000000000000001100100",
"10110010111000000000000001101010",
"10110010111000000000000001110000",
"10110010111000000000000001110110",
"10110010111000000000000001111100",
"10110010111000000000000010000010",
"10110010111000000000000010001000",
"10110010111000000000000010001110",
"11010000110000000000000000000001",
"11001000000000000000000010100110",
"10110100100000000000000010010001",
"10110100100000000000000010010100",
"01010100000100000000000000110010",
"01010100000100001000000000110010",
"10110100000000000000000010010000",
"10110100001000000000000010010011",
"11010100000000000000001111101000",
"11001000000000000000000010101001",
"11000000000000110000000000000000",
"11010000111000000000000000000001",
"11001000000000000000000010110001",
"10110100101000000000000010010111",
"10110100101000000000000010011010",
"01011100010100010000000000110010",
"01011100010100011000000000110010",
"10110100010000000000000010010110",
"10110100011000000000000010011001",
"11010100010000000111110000011000",
"11001000000000000000000010110100",
x"F0000000",
x"F0000000",
x"F0000000",
x"F0A000B0",
x"F0000000",
"11010000110000000000000000000001",
"11001000000000000000000011000001",
"11100010100000000000000000100100",
"11001000000000000000000011000001",
"11100100100000000000000000010101",
"11001000000000000000000011000001",
"11100100000000000000000000010000",
"11001000000000000000000011000001",
"11001000000000000000000011000000",
x"F0000000",
x"F0000000",
x"F0010000",
x"F0101000",
x"F0000000",
x"F0A000B0",
x"F0000000",
x"FC000000",
x"F0000000",
x"F0000000",
x"F0010000",
x"F0101000",
x"F0000000",
x"F0A000B0",
x"F0000000",
x"FC000000",
x"F0000000",
x"F0000000",
x"F0010000",
x"F0101000",
x"F0000000",
x"F0A000B0",
x"F0000000",
x"FC000000",
x"F0000000",
x"F0000000",
x"F0010000",
x"F0101000",
x"F0000000",
x"F0A000B0",
x"F0000000",
x"FC000000",
x"F0000000",
x"F0000000",
x"F0010000",
x"F0101000",
x"F0000000",
x"F0A000B0",
x"F0000000",
x"FC000000",
x"F0000000",
x"F0000000",
x"F0010000",
x"F0101000",
x"F0000000",
x"F0A000B0",
x"F0000000",
x"FC000000",
x"F0000000",
x"F0000000",
x"F0010000",
x"F0101000",
x"F0000000",
x"F0A000B0",
x"F0000000",
x"FC000000",
x"F0000000",
x"F0000000",
x"F0010000",
x"F0101000",
x"F0000000",
x"F0A000B0",
x"F0000000");

begin

process(order)begin

inst<=reg(to_integer(unsigned(order)));

end process;

end Behavioral;
